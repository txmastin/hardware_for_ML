*------------------------------------------------------------
* test_orig_memC.cir — Standalone test of Biolek memcapacitor
*------------------------------------------------------------
.option method=gear reltol=1e-4 abstol=1e-12 vntol=1e-6

* Slow sine drive (1 Hz, 2 V amplitude)
Vtest plus 0 SIN(0 2 1)

* Instantiate the memC_orig subcircuit
Xmem plus minus memC_orig Cmin=10n Cmax=10u Cinit=100n k=10meg p=1 IC=0

* Prevent floating internal nodes
Rshunt minus 0 1G
Rst_q   charge 0 1G
Rst_x   x      0 1G

* Transient run for hysteresis to develop
.tran 1ms 200ms uic

.control
  run
  * Plot terminal voltages and internal state
  plot V(plus) V(minus) V(x) V(charge)
.endc

*------------------------------------------------------------
* Original Biolek et al. 2010 memcapacitor subcircuit
*------------------------------------------------------------
.SUBCKT memC_orig plus minus Cmin=10n Cmax=10u Cinit=100n k=10meg p=1 IC=0
  * Controlled voltage: Emc = DM(x)*(q + IC·Cinit)
  Emc plus minus VALUE = { DM(V(x)) * ( V(charge) + IC * Cinit ) }

  * Charge integrator (Int1)
  Gq  0 charge VALUE = { I(Emc) }
  Cq  charge 0 1
  Rq  charge 0 1G

  * State integrator (Int2)
  .PARAM xinit = { (1/Cinit - 1/Cmax) / (1/Cmin - 1/Cmax) }
  Gx  0 x VALUE = { V(charge) * k * window(V(x), p) }
  Cx  x 0 1 IC = { xinit }
  Rx  x 0 1G

  * Core functions
  .FUNC DM(x)     = { 1/Cmax + (1/Cmin - 1/Cmax) * x }
  .FUNC window(x,p) = { 1 - pow(2*x - 1, 2*p) }
.ENDS memC_orig

