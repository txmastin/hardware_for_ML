*------------------------------------------------------------
* FLIF Neuron with Enhanced Memcapacitor
* Based on Vazquez-Guerrero (2024) + your Biolek-style memC
*------------------------------------------------------------

* Parameters
.param Vthresh = 1.5
.param Rleak = 10Meg
.param Vdd = 5

* Power supply for spike path
Vdd_node Vdd 0 DC {Vdd}

* Input current (synaptic current pulse)
Iin in 0 PULSE(0 10u 1ms 1ms 1ms 5ms 100ms)
Rin in vmem 1Meg

* Leak resistor
Rleak vmem 0 {Rleak}

* Memcapacitor (hysteretic, nonlinear)
Xmem vmem 0 memcapacitor params: Cmin=1p Cmax=10n beta=0.2 x0=0.1 p=10

* Threshold reference
Vth vthresh 0 DC {Vthresh}

* Spike detection (MOSFET-based comparator output)
* Instead of analog spike pulse, we’ll just use a behavioral spike output for now
Bspike spike_out 0 V = '10 * exp(-((V(vmem) - V(vthresh))^2) / 0.001)'

*------------------------------------------------------------
* Analysis
*------------------------------------------------------------
.tran 0.1ms 1000ms uic

.control
run
* Plot voltage and spike output
plot V(vmem) V(spike_out)
.endc

*------------------------------------------------------------
* Enhanced Memcapacitor Subcircuit
*------------------------------------------------------------
.subckt memcapacitor plus minus params:
+ Cmin=1p
+ Cmax=10n
+ beta=0.2
+ x0=0.1
+ p=10

.nodeset v(xvar)={x0}
Cx xvar 0 1

* Biolek-style window function
.func biolek_win(x,i) = {1-pow(2*x-1,2*p) * ((i>0) * (x>0.98) + (i<=0) * (x<0.02))}

* State variable evolution
Bx 0 xvar I={beta*V(plus,minus)*V(plus,minus)*biolek_win(V(xvar),V(plus,minus))}

* Capacitance as function of x
Ec cap 0 value={Cmin+((Cmax-Cmin)*pow(V(xvar),2))}

* Memcapacitive current
Gmem plus minus value={V(cap)*ddt(V(plus,minus)) + (2*(Cmax-Cmin)*V(xvar))*V(plus,minus)*I(Cx)}

.ends memcapacitor

