* Purely Hardware-Analog Leaky Integrate-and-Fire (LIF) Neuron
* Corrected resistor values for Hardware Schmitt Trigger.
* Added .NODESET directives to guide initial DC solution.

*******************************************************************************
* Parameters
*******************************************************************************
.param R_LK = 10k      ; Leak resistance (Ohms)
.param C_MEM = 100n     ; Membrane capacitance (Farads)
.param V_RESET_VAL = 0.0  ; Reset voltage value (Volts) - Vm is pulled towards this

* Op-Amp Core Parameters (for the op-amp used in Schmitt trigger)
.param VCC_OPAMP = 5.0  ; Positive rail for op-amp (Volts)
.param VEE_OPAMP = 0.0  ; Negative rail for op-amp (Volts)
.param OPAMP_GAIN_CORE = 100Meg ; Gain for the op-amp core

* Schmitt Trigger Resistor and Reference Voltage Parameters
* Designed for UTP = 1.0V, LTP = 0.2V
.param R_SCHMITT_1_PARAM = 1.6k   ; << CORRECTED: Resistor from Vm to op-amp V+
.param R_SCHMITT_2_PARAM = 10k    ; << CORRECTED: Resistor from Vcomp_out (op-amp output) to op-amp V+
.param V_REF_SCHMITT_PARAM = 0.86207 ; Reference voltage for op-amp V- (approx 1.0/1.16)

* MOSFET Parameters
.param MOSFET_VTO = 0.5  ; MOSFET Threshold Voltage (ensure 0V < VTO < 5V)
.param MOSFET_KP = 1m   ; MOSFET Transconductance (1000u)
.param MOSFET_W = 20u   ; MOSFET Width
.param MOSFET_L = 1u    ; MOSFET Length

* Input current - CONSTANT DC
.param I_CONST_IN = 190u ; Constant input current (Amps)

* Simulation parameters
.param T_STOP = 50m     ; Total simulation time
.param T_STEP = 0.1u    ; Maximum timestep (kept small)

*******************************************************************************
* Circuit Netlist
*******************************************************************************

* --- Input Current Source (Constant DC) ---
Iin 0 Vm DC {I_CONST_IN}

* --- Leaky Integrator Core ---
Rleak Vm 0 {R_LK}
Cmem  Vm 0 {C_MEM} IC={V_RESET_VAL} ; Initial condition

* --- Voltage Reference for Reset Target ---
Vreset_target_node reset_target 0 DC {V_RESET_VAL}

* --- Schmitt Trigger Circuit Components ---
* Reference voltage for the Schmitt trigger's op-amp
V_REF_SRC V_REF_SCHMITT_NODE 0 DC {V_REF_SCHMITT_PARAM}

* Resistors for Schmitt trigger positive feedback
R_SCHMITT_1 Vm Vplus_opamp_node {R_SCHMITT_1_PARAM}
R_SCHMITT_2 Vcomp_out Vplus_opamp_node {R_SCHMITT_2_PARAM}

* Op-Amp Core for Schmitt Trigger (Behavioral Model of an Op-Amp IC)
* Non-inverting input is Vplus_opamp_node, Inverting input is V_REF_SCHMITT_NODE
B_OPAMP_CORE Vcomp_out 0 V = min({VCC_OPAMP}, max({VEE_OPAMP}, {OPAMP_GAIN_CORE}*(V(Vplus_opamp_node) - V(V_REF_SCHMITT_NODE))))

* --- MOSFET Reset Switch ---
* Drain connected to Vm, Source connected to reset_target_node
* Gate driven by the output of the Schmitt trigger (Vcomp_out)
Mreset Vm Vcomp_out reset_target reset_target NMOS_RESET L={MOSFET_L} W={MOSFET_W}
.model NMOS_RESET NMOS (LEVEL=1 VTO={MOSFET_VTO} KP={MOSFET_KP} GAMMA=0.3 PHI=0.6 LAMBDA=0)

* --- Initial Condition Guidance ---
.NODESET V(Vm)={V_RESET_VAL} V(Vcomp_out)={VEE_OPAMP} V(Vplus_opamp_node)=0

*******************************************************************************
* Analysis
*******************************************************************************
.TRAN {T_STEP} {T_STOP} UIC

*******************************************************************************
* Control Block for ngspice
*******************************************************************************
.control
    run
    set NOPTS
    set noaskquit
    set color0=white
    set color1=black
    set xgridwidth=2

    plot V(Vm) title 'Membrane Potential (Corrected HW Schmitt Trigger LIF)' ylimit -0.1 1.1
    plot V(Vcomp_out) title 'Corrected HW Schmitt Trigger Output' ylimit -0.1 5.1
    plot I(Iin) title 'Input Current'
.endc

.end

