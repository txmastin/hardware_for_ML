* flif_oustaloup_final.cir — Fractional LIF via Oustaloup in NGSpice

*—— Solver Settings ——————————————————————————————
.options METHOD=GEAR RELTOL=1e-4 VNTOL=1e-6 ABSTOL=1e-12 ITL4=200

*—— Parameters —————————————————————————————————————
.param Iin_amp  = 2e-6     ; input current (A)
.param Vth      = 0.5      ; spike threshold (V)
.param Ireset   = 50e-6    ; reset current amplitude (A)

* Oustaloup coefficients for H(s)=1/(τ s^α + 1), α=0.8, N=5
.param num0=1.00000000e+00 num1=8.78886950e+03 num2=7.02157046e+06
.param num3=5.55410552e+08 num4=4.34983337e+09 num5=3.09670148e+09

.param den0=1.00050000e+00 den1=8.81659651e+03 den2=7.16133734e+06
.param den3=6.25166964e+08 den4=7.79684402e+09 den5=1.85802089e+10

*—— Circuit ——————————————————————————————————————
* 1) Convert Iin → V(dummy) via 1Ω resistor
Iin    dummy 0 DC {Iin_amp}
Rdm    dummy 0 1

* 2) Fractional membrane voltage via behavioral Laplace
*    use curly braces for coefficient lists!
Bfrac  membrane 0 V=laplace(V(dummy), {num0 num1 num2 num3 num4 num5}, {den0 den1 den2 den3 den4 den5})

* 3) Threshold reference
Vthref vth_ref 0 DC {Vth}

* 4) Comparator → control node
Bcomp   ctrl    0 V={ V(membrane)>V(vth_ref) ? 1 : 0 }
Rg      ctrl    0 1e12

* 5) Reset‐pulse current
Breset  membrane 0 I={ -Ireset * (V(ctrl)>0.5 ? 1 : 0) }

* 6) Initial conditions & simulate
.ic V(membrane)=0 V(ctrl)=0

.tran 1e-7 1e-2 uic

.control
  run
  plot V(membrane) V(ctrl) I(Breset)*1e6
.endc

.end

