* Memcapacitor Model for NGSPICE - Simplified Version
* Simple voltage-controlled memcapacitor model compatible with NGSPICE

.subckt memcapacitor plus minus params:
+ Cmin=1p      ; Minimum capacitance value (F)
+ Cmax=500p    ; Maximum capacitance value (F) - increased for more visible hysteresis
+ beta=0.05    ; Rate of change for state variable - increased for faster evolution
+ x0=0.5       ; Initial value of state variable (between 0 and 1)

* Internal node for state variable
.nodeset v(xvar)={x0}
Cx xvar 0 1

* Simpler window function implementation
.func w_up(x) = {1-(x-0.98)*(x>0.98)}
.func w_dn(x) = {1-(0.02-x)*(x<0.02)}
.func win(x,v) = {(v>0)*w_up(x) + (v<=0)*w_dn(x)}

* State variable evolution - controlled by voltage
Bx 0 xvar I={beta*V(plus,minus)*win(V(xvar),V(plus,minus))}

* Memcapacitor current implementation
Ec cap 0 value={Cmin+(Cmax-Cmin)*V(xvar)}
Gmem plus minus value={V(cap)*ddt(V(plus,minus)) + (Cmax-Cmin)*V(plus,minus)*I(Cx)}

.ends memcapacitor

* Test circuit
vsrc in 0 SIN(0 2 100)   ; 2V amplitude, 100Hz sine wave
xmem in 0 memcapacitor params: Cmin=1p Cmax=100p beta=1e-2 x0=0.5

* Analysis commands
.control
tran 0.1m 50m uic  ; Use initial conditions
let cap_state = v(xmem.xvar)   ; Save state variable
let current = i(vsrc)          ; Save current
let voltage = v(in)            ; Save voltage

* Run multiple cycles to allow state to evolve
plot voltage current*1e9       ; Plot voltage and current vs time
plot voltage vs current*1e9 retraceplot    ; Plot I-V curve to see hysteresis

* Plot multiple cycles to see evolution of hysteresis
set curplottitle="I-V Hysteresis Curve of Memcapacitor"
plot current*1e9 vs voltage xlimit -2 2 ylimit -20 20 retraceplot
.endc

.end
