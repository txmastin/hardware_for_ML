*------------------------------------------------------------
* FLIF Neuron with Enhanced Memcapacitor — Stable Version
*------------------------------------------------------------

* Global parameters
.param Vthresh = 1.5
.param Rleak   = 10Meg
.param Vdd     = 5

* Power supply for any MOSFET paths (unused here)
Vdd_node Vdd 0 DC {Vdd}

* Synaptic input: 10 µA pulse
Iin    in    0 PULSE(0 10u 100ms 1ms 1ms 200ms 1000ms)
Rin    in    vmem 1Meg

* Leak path
Rleak  vmem  0    {Rleak}

* Replace classical Cm with your enhanced memcapacitor
Xmem   vmem  0    memcapacitor params: Cmin=1p Cmax=100p beta=1e-3 x0=0.1 p=10

* Threshold reference
Vth    vth   0    DC {Vthresh}

* Behavioral spike output (Gaussian around threshold)
Bspike spike_out 0 V = '10 * exp(-((V(vmem)-V(vth))**2) / 0.001)'

* Transient and numerical settings
.tran 0.01ms 1000ms uic
.options maxstep=0.1ms

.control
  run
  plot V(vmem) V(spike_out)
.endc

*------------------------------------------------------------
* Enhanced Memcapacitor Subcircuit (stable Gmem)
*------------------------------------------------------------
.subckt memcapacitor plus minus params:
+ Cmin=1p Cmax=100p beta=1e-3 x0=0.1 p=10

* Initialize internal state xvar
.nodeset v(xvar)={x0}
Cx       xvar 0 1

* Soft clamp: xvar_limited ∈ [0,1]
Bxlim    xvar_limited 0 V = 'min(max(V(xvar),0),1)'

* Biolek directional window
.func biolek_win(x,i) = {1 - pow(2*x-1,2*p) * ((i>0)*(x>0.98) + (i<=0)*(x<0.02))}

* State evolution
Bx       0 xvar I = {beta * V(plus,minus)**2 * biolek_win(V(xvar_limited),V(plus,minus))}

* Effective capacitance node
Ec       cap 0 value = {Cmin + (Cmax - Cmin) * V(xvar_limited)**2}

* Memcapacitive current (stable)
Gmem     plus minus value = { V(cap) * ddt(V(plus,minus)) }

.ends memcapacitor

