*------------------------------------------------------------
* FLIF neuron with Biolek memcapacitor (fixed instantiation)
*------------------------------------------------------------

.param Vth    = 1.0
.param Iin_amp= 2u
.param Rin    = 1Meg
.param Rleak  = 500k
.param Ireset = 50u
.param dt     = 0.01ms
.param Tstop  = 200ms

Iin   0   in    DC {Iin_amp}
Rin   in  vmem  {Rin}
Rleak vmem 0    {Rleak}

* Correct instantiation of memcapacitor
Xmem  vmem 0   memcapacitor Cmin=10n Cmax=10u Cinit=100n k=10meg p=1 IC=0

* Fire when vmem > Vth (since you flipped it back to positive domain)
Bfire fire 0 V = 'V(vmem) > {Vth} ? 1 : 0'

* RESET as a continuous current sink
Greset vmem 0 VALUE = { V(fire) * Ireset }

Bspike spike_out 0 V = 'V(fire)*10'

.option method=gear
.option numdgt=12 reltol=1e-4 abstol=1e-9 vntol=1e-6
.tran {dt} {Tstop} uic

.control
  run
  plot V(vmem) V(spike_out)
.endc

*------------------------------------------------------------
* Biolek et al. 2010 Memcapacitor Subcircuit (renamed)
*------------------------------------------------------------
.SUBCKT memcapacitor plus minus Cmin=10n Cmax=10u Cinit=100n k=10meg p=1 IC=0
Emc plus minus VALUE={DM(V(x))*(V(charge)+IC*Cinit)}
Gq 0 charge VALUE={I(Emc)}
Cq charge 0 1
Rq charge 0 1G
.PARAM xinit={(1/Cinit-1/Cmax)/(1/Cmin-1/Cmax)}
Gx 0 x VALUE={V(charge)*k*window(V(x),p)}
Cx x 0 1 IC={xinit}
Rx x 0 1G
.FUNC DM(x)      ={1/Cmax + (1/Cmin-1/Cmax)*x}
.FUNC window(x,p)={1 - pow(2*x-1,2*p)}
.ENDS memcapacitor

